`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    07:52:14 09/06/2023 
// Design Name: 
// Module Name:    counter4bit 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module counter4bit(
    input wire clk,
    input wire reset,
    output wire [3:0] q
    );
// signal declaration
reg [3:0] r_reg;
wire [3:0] r_next;
// body, register
always @(posedge clk, posedge reset)
if (reset)
r_reg <= 0;
 else
r_reg<=r_next; // <= is non-blocking statement
// next state logic
assign r_next = r_reg + 1;
// output logic
assign q=r_reg;
endmodule



